library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
library UNISIM;
use UNISIM.VComponents.all;

entity deney4vhdl22 is
    Port ( A : in  STD_LOGIC_VECTOR (0 downto 3);
           S : out  STD_LOGIC_VECTOR (0 downto 7));
end deney4vhdl22;

architecture Behavioral of deney4vhdl22 is

begin


end Behavioral;

